----------------------------------------------------------------------------------------------------
-- Copyright (c) 2018 Marcus Geelnard
--
-- This software is provided 'as-is', without any express or implied warranty. In no event will the
-- authors be held liable for any damages arising from the use of this software.
--
-- Permission is granted to anyone to use this software for any purpose, including commercial
-- applications, and to alter it and redistribute it freely, subject to the following restrictions:
--
--  1. The origin of this software must not be misrepresented; you must not claim that you wrote
--     the original software. If you use this software in a product, an acknowledgment in the
--     product documentation would be appreciated but is not required.
--
--  2. Altered source versions must be plainly marked as such, and must not be misrepresented as
--     being the original software.
--
--  3. This notice may not be removed or altered from any source distribution.
----------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use work.common.all;

entity shift32_tb is
end shift32_tb;

architecture behavioral of shift32_tb is
  signal s_right       : std_logic;
  signal s_arithmetic  : std_logic;
  signal s_src         : std_logic_vector(31 downto 0);
  signal s_shift       : std_logic_vector(31 downto 0);
  signal s_packed_mode : T_PACKED_MODE;
  signal s_result      : std_logic_vector(31 downto 0);

  signal s_op : std_logic_vector(1 downto 0);

  function shft32(a: integer) return std_logic_vector is
  begin
    return to_vector(a, 32);
  end function;

  function shft16(a: integer; b: integer) return std_logic_vector is
  begin
    return to_vector(a, 16) & to_vector(b, 16);
  end function;

  function shft8(a: integer; b: integer; c: integer; d: integer) return std_logic_vector is
  begin
    return to_vector(a, 8) & to_vector(b, 8) & to_vector(c, 8) & to_vector(d, 8);
  end function;

begin
  shift32_0: entity work.shift32
    port map (
      i_right => s_right,
      i_arithmetic => s_arithmetic,
      i_src => s_src,
      i_shift => s_shift,
      i_packed_mode => s_packed_mode,
      o_result => s_result
    );

  process
    --  The patterns to apply.
    type pattern_type is record
      -- Inputs
      right       : std_logic;
      arithmetic  : std_logic;
      src         : std_logic_vector(31 downto 0);
      shift       : std_logic_vector(31 downto 0);
      packed_mode : T_PACKED_MODE;

      -- Expected outputs
      result     : std_logic_vector(31 downto 0);
    end record;
    type pattern_array is array (natural range <>) of pattern_type;
    constant patterns : pattern_array := (
        -- LSL
        ('0', '0', "10001111000001110000001100000001", shft32(0), C_PACKED_NONE, "10001111000001110000001100000001"),
        ('0', '0', "10001111000001110000001100000001", shft32(1), C_PACKED_NONE, "00011110000011100000011000000010"),
        ('0', '0', "10001111000001110000001100000001", shft32(2), C_PACKED_NONE, "00111100000111000000110000000100"),
        ('0', '0', "10001111000001110000001100000001", shft32(3), C_PACKED_NONE, "01111000001110000001100000001000"),
        ('0', '0', "10001111000001110000001100000001", shft32(4), C_PACKED_NONE, "11110000011100000011000000010000"),
        ('0', '0', "10001111000001110000001100000001", shft32(5), C_PACKED_NONE, "11100000111000000110000000100000"),
        ('0', '0', "10001111000001110000001100000001", shft32(6), C_PACKED_NONE, "11000001110000001100000001000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(7), C_PACKED_NONE, "10000011100000011000000010000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(8), C_PACKED_NONE, "00000111000000110000000100000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(9), C_PACKED_NONE, "00001110000001100000001000000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(10), C_PACKED_NONE, "00011100000011000000010000000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(11), C_PACKED_NONE, "00111000000110000000100000000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(12), C_PACKED_NONE, "01110000001100000001000000000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(13), C_PACKED_NONE, "11100000011000000010000000000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(14), C_PACKED_NONE, "11000000110000000100000000000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(15), C_PACKED_NONE, "10000001100000001000000000000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(16), C_PACKED_NONE, "00000011000000010000000000000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(17), C_PACKED_NONE, "00000110000000100000000000000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(18), C_PACKED_NONE, "00001100000001000000000000000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(19), C_PACKED_NONE, "00011000000010000000000000000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(20), C_PACKED_NONE, "00110000000100000000000000000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(21), C_PACKED_NONE, "01100000001000000000000000000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(22), C_PACKED_NONE, "11000000010000000000000000000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(23), C_PACKED_NONE, "10000000100000000000000000000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(24), C_PACKED_NONE, "00000001000000000000000000000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(25), C_PACKED_NONE, "00000010000000000000000000000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(26), C_PACKED_NONE, "00000100000000000000000000000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(27), C_PACKED_NONE, "00001000000000000000000000000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(28), C_PACKED_NONE, "00010000000000000000000000000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(29), C_PACKED_NONE, "00100000000000000000000000000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(30), C_PACKED_NONE, "01000000000000000000000000000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(31), C_PACKED_NONE, "10000000000000000000000000000000"),
        ('0', '0', "10001111000001110000001100000001", shft32(32), C_PACKED_NONE, "10001111000001110000001100000001"),
        ('0', '0', "10001111000001110000001100000001", shft32(33), C_PACKED_NONE, "00011110000011100000011000000010"),

        ('0', '0', "10001111000001111000001100000001", shft16(0, 1), C_PACKED_HALF_WORD, "10001111000001110000011000000010"),
        ('0', '0', "10001111000001111000001100000001", shft16(2, 3), C_PACKED_HALF_WORD, "00111100000111000001100000001000"),
        ('0', '0', "10001111000001111000001100000001", shft16(4, 5), C_PACKED_HALF_WORD, "11110000011100000110000000100000"),
        ('0', '0', "10001111000001111000001100000001", shft16(6, 7), C_PACKED_HALF_WORD, "11000001110000001000000010000000"),
        ('0', '0', "10001111000001111000001100000001", shft16(8, 9), C_PACKED_HALF_WORD, "00000111000000000000001000000000"),
        ('0', '0', "10001111000001111000001100000001", shft16(10, 11), C_PACKED_HALF_WORD, "00011100000000000000100000000000"),
        ('0', '0', "10001111000001111000001100000001", shft16(12, 13), C_PACKED_HALF_WORD, "01110000000000000010000000000000"),
        ('0', '0', "10001111000001111000001100000001", shft16(14, 15), C_PACKED_HALF_WORD, "11000000000000001000000000000000"),
        ('0', '0', "10001111000001111000001100000001", shft16(16, 17), C_PACKED_HALF_WORD, "10001111000001110000011000000010"),

        ('0', '0', "10001111100001111000001110000001", shft8(0, 1, 2, 3), C_PACKED_BYTE, "10001111000011100000110000001000"),
        ('0', '0', "10001111100001111000001110000001", shft8(4, 5, 6, 7), C_PACKED_BYTE, "11110000111000001100000010000000"),
        ('0', '0', "10001111100001111000001110000001", shft8(8, 9, 10, 11), C_PACKED_BYTE, "10001111000011100000110000001000"),

        -- LSR
        ('1', '0', "10001111000001110000001100000001", shft32(0), C_PACKED_NONE, "10001111000001110000001100000001"),
        ('1', '0', "10001111000001110000001100000001", shft32(1), C_PACKED_NONE, "01000111100000111000000110000000"),
        ('1', '0', "10001111000001110000001100000001", shft32(2), C_PACKED_NONE, "00100011110000011100000011000000"),
        ('1', '0', "10001111000001110000001100000001", shft32(3), C_PACKED_NONE, "00010001111000001110000001100000"),
        ('1', '0', "10001111000001110000001100000001", shft32(4), C_PACKED_NONE, "00001000111100000111000000110000"),
        ('1', '0', "10001111000001110000001100000001", shft32(5), C_PACKED_NONE, "00000100011110000011100000011000"),
        ('1', '0', "10001111000001110000001100000001", shft32(6), C_PACKED_NONE, "00000010001111000001110000001100"),
        ('1', '0', "10001111000001110000001100000001", shft32(7), C_PACKED_NONE, "00000001000111100000111000000110"),
        ('1', '0', "10001111000001110000001100000001", shft32(8), C_PACKED_NONE, "00000000100011110000011100000011"),
        ('1', '0', "10001111000001110000001100000001", shft32(9), C_PACKED_NONE, "00000000010001111000001110000001"),
        ('1', '0', "10001111000001110000001100000001", shft32(10), C_PACKED_NONE, "00000000001000111100000111000000"),
        ('1', '0', "10001111000001110000001100000001", shft32(11), C_PACKED_NONE, "00000000000100011110000011100000"),
        ('1', '0', "10001111000001110000001100000001", shft32(12), C_PACKED_NONE, "00000000000010001111000001110000"),
        ('1', '0', "10001111000001110000001100000001", shft32(13), C_PACKED_NONE, "00000000000001000111100000111000"),
        ('1', '0', "10001111000001110000001100000001", shft32(14), C_PACKED_NONE, "00000000000000100011110000011100"),
        ('1', '0', "10001111000001110000001100000001", shft32(15), C_PACKED_NONE, "00000000000000010001111000001110"),
        ('1', '0', "10001111000001110000001100000001", shft32(16), C_PACKED_NONE, "00000000000000001000111100000111"),
        ('1', '0', "10001111000001110000001100000001", shft32(17), C_PACKED_NONE, "00000000000000000100011110000011"),
        ('1', '0', "10001111000001110000001100000001", shft32(18), C_PACKED_NONE, "00000000000000000010001111000001"),
        ('1', '0', "10001111000001110000001100000001", shft32(19), C_PACKED_NONE, "00000000000000000001000111100000"),
        ('1', '0', "10001111000001110000001100000001", shft32(20), C_PACKED_NONE, "00000000000000000000100011110000"),
        ('1', '0', "10001111000001110000001100000001", shft32(21), C_PACKED_NONE, "00000000000000000000010001111000"),
        ('1', '0', "10001111000001110000001100000001", shft32(22), C_PACKED_NONE, "00000000000000000000001000111100"),
        ('1', '0', "10001111000001110000001100000001", shft32(23), C_PACKED_NONE, "00000000000000000000000100011110"),
        ('1', '0', "10001111000001110000001100000001", shft32(24), C_PACKED_NONE, "00000000000000000000000010001111"),
        ('1', '0', "10001111000001110000001100000001", shft32(25), C_PACKED_NONE, "00000000000000000000000001000111"),
        ('1', '0', "10001111000001110000001100000001", shft32(26), C_PACKED_NONE, "00000000000000000000000000100011"),
        ('1', '0', "10001111000001110000001100000001", shft32(27), C_PACKED_NONE, "00000000000000000000000000010001"),
        ('1', '0', "10001111000001110000001100000001", shft32(28), C_PACKED_NONE, "00000000000000000000000000001000"),
        ('1', '0', "10001111000001110000001100000001", shft32(29), C_PACKED_NONE, "00000000000000000000000000000100"),
        ('1', '0', "10001111000001110000001100000001", shft32(30), C_PACKED_NONE, "00000000000000000000000000000010"),
        ('1', '0', "10001111000001110000001100000001", shft32(31), C_PACKED_NONE, "00000000000000000000000000000001"),
        ('1', '0', "10001111000001110000001100000001", shft32(32), C_PACKED_NONE, "10001111000001110000001100000001"),
        ('1', '0', "10001111000001110000001100000001", shft32(33), C_PACKED_NONE, "01000111100000111000000110000000"),

        ('1', '0', "10001111000001111000001100000001", shft16(0, 1), C_PACKED_HALF_WORD, "10001111000001110100000110000000"),
        ('1', '0', "10001111000001111000001100000001", shft16(2, 3), C_PACKED_HALF_WORD, "00100011110000010001000001100000"),
        ('1', '0', "10001111000001111000001100000001", shft16(4, 5), C_PACKED_HALF_WORD, "00001000111100000000010000011000"),
        ('1', '0', "10001111000001111000001100000001", shft16(6, 7), C_PACKED_HALF_WORD, "00000010001111000000000100000110"),
        ('1', '0', "10001111000001111000001100000001", shft16(8, 9), C_PACKED_HALF_WORD, "00000000100011110000000001000001"),
        ('1', '0', "10001111000001111000001100000001", shft16(10, 11), C_PACKED_HALF_WORD, "00000000001000110000000000010000"),
        ('1', '0', "10001111000001111000001100000001", shft16(12, 13), C_PACKED_HALF_WORD, "00000000000010000000000000000100"),
        ('1', '0', "10001111000001111000001100000001", shft16(14, 15), C_PACKED_HALF_WORD, "00000000000000100000000000000001"),
        ('1', '0', "10001111000001111000001100000001", shft16(16, 17), C_PACKED_HALF_WORD, "10001111000001110100000110000000"),

        ('1', '0', "10001111100001111000001110000001", shft8(0, 1, 2, 3), C_PACKED_BYTE, "10001111010000110010000000010000"),
        ('1', '0', "10001111100001111000001110000001", shft8(4, 5, 6, 7), C_PACKED_BYTE, "00001000000001000000001000000001"),
        ('1', '0', "10001111100001111000001110000001", shft8(8, 9, 10, 11), C_PACKED_BYTE, "10001111010000110010000000010000"),

        -- ASR
        ('1', '1', "10001111000001110000001100000001", shft32(0), C_PACKED_NONE, "10001111000001110000001100000001"),
        ('1', '1', "10001111000001110000001100000001", shft32(1), C_PACKED_NONE, "11000111100000111000000110000000"),
        ('1', '1', "10001111000001110000001100000001", shft32(2), C_PACKED_NONE, "11100011110000011100000011000000"),
        ('1', '1', "10001111000001110000001100000001", shft32(3), C_PACKED_NONE, "11110001111000001110000001100000"),
        ('1', '1', "10001111000001110000001100000001", shft32(4), C_PACKED_NONE, "11111000111100000111000000110000"),
        ('1', '1', "10001111000001110000001100000001", shft32(5), C_PACKED_NONE, "11111100011110000011100000011000"),
        ('1', '1', "10001111000001110000001100000001", shft32(6), C_PACKED_NONE, "11111110001111000001110000001100"),
        ('1', '1', "10001111000001110000001100000001", shft32(7), C_PACKED_NONE, "11111111000111100000111000000110"),
        ('1', '1', "10001111000001110000001100000001", shft32(8), C_PACKED_NONE, "11111111100011110000011100000011"),
        ('1', '1', "10001111000001110000001100000001", shft32(9), C_PACKED_NONE, "11111111110001111000001110000001"),
        ('1', '1', "10001111000001110000001100000001", shft32(10), C_PACKED_NONE, "11111111111000111100000111000000"),
        ('1', '1', "10001111000001110000001100000001", shft32(11), C_PACKED_NONE, "11111111111100011110000011100000"),
        ('1', '1', "10001111000001110000001100000001", shft32(12), C_PACKED_NONE, "11111111111110001111000001110000"),
        ('1', '1', "10001111000001110000001100000001", shft32(13), C_PACKED_NONE, "11111111111111000111100000111000"),
        ('1', '1', "10001111000001110000001100000001", shft32(14), C_PACKED_NONE, "11111111111111100011110000011100"),
        ('1', '1', "10001111000001110000001100000001", shft32(15), C_PACKED_NONE, "11111111111111110001111000001110"),
        ('1', '1', "10001111000001110000001100000001", shft32(16), C_PACKED_NONE, "11111111111111111000111100000111"),
        ('1', '1', "10001111000001110000001100000001", shft32(17), C_PACKED_NONE, "11111111111111111100011110000011"),
        ('1', '1', "10001111000001110000001100000001", shft32(18), C_PACKED_NONE, "11111111111111111110001111000001"),
        ('1', '1', "10001111000001110000001100000001", shft32(19), C_PACKED_NONE, "11111111111111111111000111100000"),
        ('1', '1', "10001111000001110000001100000001", shft32(20), C_PACKED_NONE, "11111111111111111111100011110000"),
        ('1', '1', "10001111000001110000001100000001", shft32(21), C_PACKED_NONE, "11111111111111111111110001111000"),
        ('1', '1', "10001111000001110000001100000001", shft32(22), C_PACKED_NONE, "11111111111111111111111000111100"),
        ('1', '1', "10001111000001110000001100000001", shft32(23), C_PACKED_NONE, "11111111111111111111111100011110"),
        ('1', '1', "10001111000001110000001100000001", shft32(24), C_PACKED_NONE, "11111111111111111111111110001111"),
        ('1', '1', "10001111000001110000001100000001", shft32(25), C_PACKED_NONE, "11111111111111111111111111000111"),
        ('1', '1', "10001111000001110000001100000001", shft32(26), C_PACKED_NONE, "11111111111111111111111111100011"),
        ('1', '1', "10001111000001110000001100000001", shft32(27), C_PACKED_NONE, "11111111111111111111111111110001"),
        ('1', '1', "10001111000001110000001100000001", shft32(28), C_PACKED_NONE, "11111111111111111111111111111000"),
        ('1', '1', "10001111000001110000001100000001", shft32(29), C_PACKED_NONE, "11111111111111111111111111111100"),
        ('1', '1', "10001111000001110000001100000001", shft32(30), C_PACKED_NONE, "11111111111111111111111111111110"),
        ('1', '1', "10001111000001110000001100000001", shft32(31), C_PACKED_NONE, "11111111111111111111111111111111"),
        ('1', '1', "10001111000001110000001100000001", shft32(32), C_PACKED_NONE, "10001111000001110000001100000001"),
        ('1', '1', "10001111000001110000001100000001", shft32(33), C_PACKED_NONE, "11000111100000111000000110000000"),

        ('1', '1', "10001111000001111000001100000001", shft16(0, 1), C_PACKED_HALF_WORD, "10001111000001111100000110000000"),
        ('1', '1', "10001111000001111000001100000001", shft16(2, 3), C_PACKED_HALF_WORD, "11100011110000011111000001100000"),
        ('1', '1', "10001111000001111000001100000001", shft16(4, 5), C_PACKED_HALF_WORD, "11111000111100001111110000011000"),
        ('1', '1', "10001111000001111000001100000001", shft16(6, 7), C_PACKED_HALF_WORD, "11111110001111001111111100000110"),
        ('1', '1', "10001111000001111000001100000001", shft16(8, 9), C_PACKED_HALF_WORD, "11111111100011111111111111000001"),
        ('1', '1', "10001111000001111000001100000001", shft16(10, 11), C_PACKED_HALF_WORD, "11111111111000111111111111110000"),
        ('1', '1', "10001111000001111000001100000001", shft16(12, 13), C_PACKED_HALF_WORD, "11111111111110001111111111111100"),
        ('1', '1', "10001111000001111000001100000001", shft16(14, 15), C_PACKED_HALF_WORD, "11111111111111101111111111111111"),
        ('1', '1', "10001111000001111000001100000001", shft16(16, 17), C_PACKED_HALF_WORD, "10001111000001111100000110000000"),

        ('1', '1', "10001111100001111000001110000001", shft8(0, 1, 2, 3), C_PACKED_BYTE, "10001111110000111110000011110000"),
        ('1', '1', "10001111100001111000001110000001", shft8(4, 5, 6, 7), C_PACKED_BYTE, "11111000111111001111111011111111"),
        ('1', '1', "10001111100001111000001110000001", shft8(8, 9, 10, 11), C_PACKED_BYTE, "10001111110000111110000011110000")
      );
  begin
    -- Test all the patterns in the pattern array.
    for i in patterns'range loop
      --  Set the inputs.
      s_right <= patterns(i).right;
      s_arithmetic <= patterns(i).arithmetic;
      s_src <= patterns(i).src;
      s_shift <= patterns(i).shift;
      s_packed_mode <= patterns(i).packed_mode;

      --  Wait for the results.
      wait for 1 ns;

      --  Check the outputs.
      s_op <= s_right & s_arithmetic;
      assert s_result = patterns(i).result
        report "Bad shift result:" & lf &
               "  op=" & to_string(s_op) & " shift=" & to_string(s_shift) & " pm=" & to_string(s_packed_mode) & lf &
               "  src=" & to_string(s_src) & lf &
               "  res=" & to_string(s_result) & lf &
               " (exp=" & to_string(patterns(i).result) & ")"
          severity error;
    end loop;
    assert false report "End of test" severity note;
    --  Wait forever; this will finish the simulation.
    wait;
  end process;
end behavioral;

