----------------------------------------------------------------------------------------------------
-- Copyright (c) 2018 Marcus Geelnard
--
-- This software is provided 'as-is', without any express or implied warranty. In no event will the
-- authors be held liable for any damages arising from the use of this software.
--
-- Permission is granted to anyone to use this software for any purpose, including commercial
-- applications, and to alter it and redistribute it freely, subject to the following restrictions:
--
--  1. The origin of this software must not be misrepresented; you must not claim that you wrote
--     the original software. If you use this software in a product, an acknowledgment in the
--     product documentation would be appreciated but is not required.
--
--  2. Altered source versions must be plainly marked as such, and must not be misrepresented as
--     being the original software.
--
--  3. This notice may not be removed or altered from any source distribution.
----------------------------------------------------------------------------------------------------

----------------------------------------------------------------------------------------------------
-- Pipeline Stages 4 & 5: Execute (EX1/EX2)
----------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use work.common.all;

entity execute is
  port(
    -- Control signals.
    i_clk : in std_logic;
    i_rst : in std_logic;
    o_stall : out std_logic;

    -- From ID stage (sync).
    i_pc : in std_logic_vector(C_WORD_SIZE-1 downto 0);
    i_src_a : in std_logic_vector(C_WORD_SIZE-1 downto 0);
    i_src_b : in std_logic_vector(C_WORD_SIZE-1 downto 0);
    i_src_c : in std_logic_vector(C_WORD_SIZE-1 downto 0);
    i_dst_reg : in std_logic_vector(C_LOG2_NUM_REGS-1 downto 0);
    i_writes_to_reg : in std_logic;
    i_alu_op : in T_ALU_OP;
    i_muldiv_op : in T_MULDIV_OP;
    i_mem_op : in T_MEM_OP;
    i_alu_en : in std_logic;
    i_muldiv_en : in std_logic;
    i_mem_en : in std_logic;

    -- PC signal from IF (sync).
    i_if_pc : in std_logic_vector(C_WORD_SIZE-1 downto 0);

    -- Branch signals from ID (sync).
    i_branch_reg_addr : in std_logic_vector(C_WORD_SIZE-1 downto 0);
    i_branch_offset_addr : in std_logic_vector(C_WORD_SIZE-1 downto 0);
    i_branch_is_branch : in std_logic;
    i_branch_is_reg : in std_logic;  -- 1 for register branches, 0 for all other instructions.
    i_branch_is_taken : in std_logic;

    -- Branch signals to PC (async).
    o_pccorr_target : out std_logic_vector(C_WORD_SIZE-1 downto 0);
    o_pccorr_source : out std_logic_vector(C_WORD_SIZE-1 downto 0);
    o_pccorr_is_branch : out std_logic;
    o_pccorr_is_taken : out std_logic;
    o_pccorr_adjust : out std_logic;
    o_pccorr_adjusted_pc : out std_logic_vector(C_WORD_SIZE-1 downto 0);

    -- DCache interface.
    o_dcache_req : out std_logic;  -- 1 = request, 0 = nop
    o_dcache_we : out std_logic;   -- 1 = write, 0 = read
    o_dcache_byte_mask : out std_logic_vector(C_WORD_SIZE/8-1 downto 0);
    o_dcache_addr : out std_logic_vector(C_WORD_SIZE-1 downto 2);
    o_dcache_write_data : out std_logic_vector(C_WORD_SIZE-1 downto 0);
    i_dcache_read_data : in std_logic_vector(C_WORD_SIZE-1 downto 0);
    i_dcache_read_data_ready : in std_logic;

    -- To the WB stage (sync).
    o_result : out std_logic_vector(C_WORD_SIZE-1 downto 0);
    o_dst_reg : out std_logic_vector(C_LOG2_NUM_REGS-1 downto 0);
    o_writes_to_reg : out std_logic;

    -- To operand forward logic (async).
    o_ex1_next_dst_reg : out std_logic_vector(C_LOG2_NUM_REGS-1 downto 0);
    o_ex1_next_writes_to_reg : out std_logic;
    o_ex1_next_result : out std_logic_vector(C_WORD_SIZE-1 downto 0);
    o_ex1_next_result_ready : out std_logic;
    o_ex2_next_result : out std_logic_vector(C_WORD_SIZE-1 downto 0);

    -- To operand forward logic (sync).
    o_ex1_dst_reg : out std_logic_vector(C_LOG2_NUM_REGS-1 downto 0);
    o_ex1_writes_to_reg : out std_logic;
    o_ex1_result : out std_logic_vector(C_WORD_SIZE-1 downto 0);
    o_ex1_result_ready : out std_logic
  );
end execute;

architecture rtl of execute is
  signal s_alu_result : std_logic_vector(C_WORD_SIZE-1 downto 0);

  signal s_muldiv_result : std_logic_vector(C_WORD_SIZE-1 downto 0);
  signal s_muldiv_result_ready : std_logic;
  signal s_stall_for_muldiv : std_logic;

  -- Should the EX1 stage be stalled by the EX2 stage?
  signal s_stall_ex1 : std_logic;

  -- Multicycle operation handling.
  signal s_start_multicycle_op : std_logic;
  signal s_start_muldiv_op : std_logic;
  signal s_stall_for_multicycle_op : std_logic;
  signal s_multicycle_op_finished : std_logic;
  signal s_prev_stall_for_multicycle_op : std_logic;

  signal s_next_result : std_logic_vector(C_WORD_SIZE-1 downto 0);
  signal s_next_result_ready : std_logic;

  -- Signals related to memory I/O.
  signal s_mem_byte_mask_unshifted : std_logic_vector(C_WORD_SIZE/8-1 downto 0);
  signal s_mem_byte_mask : std_logic_vector(C_WORD_SIZE/8-1 downto 0);
  signal s_mem_store_data : std_logic_vector(C_WORD_SIZE-1 downto 0);

  -- Signals for handling bubbling.
  signal s_bubble : std_logic;
  signal s_mem_op_masked : T_MEM_OP;
  signal s_mem_en_masked : std_logic;
  signal s_dst_reg_masked : std_logic_vector(C_LOG2_NUM_REGS-1 downto 0);
  signal s_writes_to_reg_masked : std_logic;

  -- Branch/PC correction signals.
  signal s_branch_target : std_logic_vector(C_WORD_SIZE-1 downto 0);
  signal s_pc_plus_4 : std_logic_vector(C_WORD_SIZE-1 downto 0);
  signal s_actual_pc : std_logic_vector(C_WORD_SIZE-1 downto 0);
  signal s_mispredicted_pc : std_logic;

  -- Signals from the EX1 to the EX2 stage (sync).
  signal s_ex1_mem_op : T_MEM_OP;
  signal s_ex1_mem_enable : std_logic;
  signal s_ex1_mem_we : std_logic;
  signal s_ex1_mem_byte_mask : std_logic_vector(C_WORD_SIZE/8-1 downto 0);
  signal s_ex1_result : std_logic_vector(C_WORD_SIZE-1 downto 0);
  signal s_ex1_result_ready : std_logic;
  signal s_ex1_store_data : std_logic_vector(C_WORD_SIZE-1 downto 0);
  signal s_ex1_dst_reg : std_logic_vector(C_LOG2_NUM_REGS-1 downto 0);
  signal s_ex1_writes_to_reg : std_logic;

  -- Signals from the memory interface (async).
  signal s_mem_stall : std_logic;
  signal s_mem_data : std_logic_vector(C_WORD_SIZE-1 downto 0);

  -- Signals from the EX2 stage (async).
  signal s_ex2_stall : std_logic;
  signal s_ex2_next_result : std_logic_vector(C_WORD_SIZE-1 downto 0);

  constant C_MULDIV_ZERO : T_MULDIV_OP := (others => '0');
begin
  --------------------------------------------------------------------------------------------------
  -- Branch logic.
  --------------------------------------------------------------------------------------------------

  -- Calculate the expected PC if no branch is taken (i.e. PC + 4).
  -- NOTE(m): We could perform this addition in the ID stage instead to save in on gate
  -- delay, at the cost of more registers.
  pc_plus_4_0: entity work.pc_plus_4
    port map (
      i_pc => i_pc,
      o_result => s_pc_plus_4
    );

  -- Check if the PC was correctly predicted by the PC stage.
  s_branch_target <= i_branch_reg_addr when i_branch_is_reg = '1' else i_branch_offset_addr;
  s_actual_pc <= s_branch_target when (i_branch_is_branch and i_branch_is_taken) = '1' else s_pc_plus_4;
  s_mispredicted_pc <= '0' when s_actual_pc = i_if_pc else i_branch_is_branch;

  -- Branch/PC correction signals to the PC stage.
  o_pccorr_target <= s_branch_target;
  o_pccorr_source <= i_pc;
  o_pccorr_is_branch <= i_branch_is_branch;
  o_pccorr_is_taken <= i_branch_is_taken;
  o_pccorr_adjust <= s_mispredicted_pc;
  o_pccorr_adjusted_pc <= s_actual_pc;


  --------------------------------------------------------------------------------------------------
  -- EX1: Execution units.
  --------------------------------------------------------------------------------------------------

  -- Should the EX1 stage be stalled?

  -- Instantiate the ALU.
  alu_1: entity work.alu
    port map (
      i_op => i_alu_op,
      i_src_a => i_src_a,
      i_src_b => i_src_b,
      o_result => s_alu_result
    );

  -- Instantiate a multiply unit.
  muldiv_1: entity work.muldiv
    port map (
      i_clk => i_clk,
      i_rst => i_rst,
      i_stall => s_stall_ex1,
      o_stall => s_stall_for_muldiv,
      i_enable => i_muldiv_en,
      i_op => i_muldiv_op,
      i_src_a => i_src_a,
      i_src_b => i_src_b,
      i_start_op => s_start_muldiv_op,
      o_result => s_muldiv_result,
      o_result_ready => s_muldiv_result_ready
    );

  -- Multicycle operation.
  s_start_multicycle_op <= i_muldiv_en and not s_prev_stall_for_multicycle_op;
  s_start_muldiv_op <= s_start_multicycle_op and i_muldiv_en;
  s_stall_for_multicycle_op <= s_stall_for_muldiv;
  s_multicycle_op_finished <= s_muldiv_result_ready;

  -- Prepare the byte mask for the MEM stage.
  ByteMaskMux: with i_mem_op(1 downto 0) select
    s_mem_byte_mask_unshifted <=
      "0001" when "01",    -- byte
      "0011" when "10",    -- halfword
      "1111" when others;  -- word (11) and undefined (00)

  ByteMaskShiftMux: with s_alu_result(1 downto 0) select
    s_mem_byte_mask <=
      s_mem_byte_mask_unshifted(3 downto 0)         when "00",
      s_mem_byte_mask_unshifted(2 downto 0) & "0"   when "01",
      s_mem_byte_mask_unshifted(1 downto 0) & "00"  when "10",
      s_mem_byte_mask_unshifted(0 downto 0) & "000" when others;  -- "11"

  -- Prepare the store data for the MEM stage (shift it into position).
  StoreDataShiftMux: with s_alu_result(1 downto 0) select
    s_mem_store_data <=
      i_src_c(31 downto 0)             when "00",
      i_src_c(23 downto 0) & X"00"     when "01",
      i_src_c(15 downto 0) & X"0000"   when "10",
      i_src_c(7 downto 0)  & X"000000" when others;  -- "11"

  -- Select the output.
  s_next_result <=
      s_alu_result when i_alu_en = '1' else
      s_muldiv_result when i_muldiv_en = '1' else
      (others => '0');

  s_next_result_ready <= (i_alu_en and (not i_mem_en)) or s_multicycle_op_finished;

  -- Should we send a bubble down the pipeline?
  -- TODO(m): We also need to bubble if there was a branch misprediction (important for not
  -- writing to LR for conditional link branches)!
  s_bubble <= s_stall_for_multicycle_op;
  s_mem_op_masked <= i_mem_op when s_bubble = '0' else (others => '0');
  s_mem_en_masked <= i_mem_en and not s_bubble;
  s_dst_reg_masked <= i_dst_reg when s_bubble = '0' else (others => '0');
  s_writes_to_reg_masked <= i_writes_to_reg and not s_bubble;

  -- Internal state.
  process(i_clk, i_rst)
  begin
    if i_rst = '1' then
      s_prev_stall_for_multicycle_op <= '0';
    elsif rising_edge(i_clk) then
      if s_stall_ex1 = '0' then
        s_prev_stall_for_multicycle_op <= s_stall_for_multicycle_op;
      end if;
    end if;
  end process;

  -- Outputs to the EX2 stage (sync).
  process(i_clk, i_rst)
  begin
    if i_rst = '1' then
      s_ex1_mem_op <= (others => '0');
      s_ex1_mem_enable <= '0';
      s_ex1_mem_we <= '0';
      s_ex1_mem_byte_mask <= (others => '0');
      s_ex1_result <= (others => '0');
      s_ex1_result_ready <= '0';
      s_ex1_store_data <= (others => '0');
      s_ex1_dst_reg <= (others => '0');
      s_ex1_writes_to_reg <= '0';
    elsif rising_edge(i_clk) then
      if s_stall_ex1 = '0' then
        s_ex1_mem_op <= s_mem_op_masked;
        s_ex1_mem_enable <= s_mem_en_masked;
        s_ex1_mem_we <= s_mem_op_masked(3);
        s_ex1_mem_byte_mask <= s_mem_byte_mask;
        s_ex1_result <= s_next_result;
        s_ex1_result_ready <= s_next_result_ready;
        s_ex1_store_data <= s_mem_store_data;
        s_ex1_dst_reg <= s_dst_reg_masked;
        s_ex1_writes_to_reg <= s_writes_to_reg_masked;
      end if;
    end if;
  end process;

  -- Output the EX1 result to operand forwarding logic.
  -- Async:
  o_ex1_next_dst_reg <= s_dst_reg_masked;
  o_ex1_next_writes_to_reg <= s_writes_to_reg_masked;
  o_ex1_next_result <= s_next_result;
  o_ex1_next_result_ready <= s_next_result_ready;

  -- Sync:
  o_ex1_dst_reg <= s_ex1_dst_reg;
  o_ex1_writes_to_reg <= s_ex1_writes_to_reg;
  o_ex1_result <= s_ex1_result;
  o_ex1_result_ready <= s_ex1_result_ready;


  --------------------------------------------------------------------------------------------------
  -- EX2: Memory.
  --------------------------------------------------------------------------------------------------

  memory_0: entity work.memory
    port map (
      o_stall => s_mem_stall,

      -- From EX1 stage (sync).
      i_mem_op => s_ex1_mem_op,
      i_mem_enable => s_ex1_mem_enable,
      i_mem_we => s_ex1_mem_we,
      i_mem_byte_mask => s_ex1_mem_byte_mask,
      i_mem_addr => s_ex1_result,
      i_store_data => s_ex1_store_data,

      -- DCache interface.
      o_dcache_req => o_dcache_req,
      o_dcache_we => o_dcache_we,
      o_dcache_byte_mask => o_dcache_byte_mask,
      o_dcache_addr => o_dcache_addr,
      o_dcache_write_data => o_dcache_write_data,
      i_dcache_read_data => i_dcache_read_data,
      i_dcache_read_data_ready => i_dcache_read_data_ready,

      -- Memory read data (async).
      o_data => s_mem_data
    );

  -- Select the result from the EX2 stage.
  s_ex2_next_result <= s_mem_data when s_ex1_mem_enable = '1' else s_ex1_result;

  -- Outputs to the WB stage (sync).
  process(i_clk, i_rst)
  begin
    if i_rst = '1' then
      o_result <= (others => '0');
      o_dst_reg <= (others => '0');
      o_writes_to_reg <= '0';
    elsif rising_edge(i_clk) then
      o_result <= s_ex2_next_result;
      o_dst_reg <= s_ex1_dst_reg;
      o_writes_to_reg <= s_ex1_writes_to_reg;
    end if;
  end process;

  -- Output the EX2 result to operand forwarding logic (async).
  o_ex2_next_result <= s_ex2_next_result;

  -- Stall logic (async).
  s_ex2_stall <= s_mem_stall;
  s_stall_ex1 <= s_ex2_stall;
  o_stall <= s_stall_for_multicycle_op or s_stall_ex1;
end rtl;

